-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80c2",
     9 => x"fc080b0b",
    10 => x"80c38008",
    11 => x"0b0b80c3",
    12 => x"84080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"c3840c0b",
    16 => x"0b80c380",
    17 => x"0c0b0b80",
    18 => x"c2fc0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbaf0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80c2fc70",
    57 => x"80cdcc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5187e3",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80c3",
    65 => x"8c0c9f0b",
    66 => x"80c3900c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"c39008ff",
    70 => x"0580c390",
    71 => x"0c80c390",
    72 => x"088025e8",
    73 => x"3880c38c",
    74 => x"08ff0580",
    75 => x"c38c0c80",
    76 => x"c38c0880",
    77 => x"25d03880",
    78 => x"0b80c390",
    79 => x"0c800b80",
    80 => x"c38c0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80c38c08",
   100 => x"25913882",
   101 => x"c82d80c3",
   102 => x"8c08ff05",
   103 => x"80c38c0c",
   104 => x"838a0480",
   105 => x"c38c0880",
   106 => x"c3900853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80c38c08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"c3900881",
   116 => x"0580c390",
   117 => x"0c80c390",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80c390",
   121 => x"0c80c38c",
   122 => x"08810580",
   123 => x"c38c0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480c3",
   128 => x"90088105",
   129 => x"80c3900c",
   130 => x"80c39008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80c390",
   134 => x"0c80c38c",
   135 => x"08810580",
   136 => x"c38c0c02",
   137 => x"8c050d04",
   138 => x"02ec050d",
   139 => x"800b80c3",
   140 => x"940cf68c",
   141 => x"08f69008",
   142 => x"71882c56",
   143 => x"5481ff06",
   144 => x"52737225",
   145 => x"89387154",
   146 => x"820b80c3",
   147 => x"940c7288",
   148 => x"2c7381ff",
   149 => x"06545574",
   150 => x"73258d38",
   151 => x"7280c394",
   152 => x"08840780",
   153 => x"c3940c55",
   154 => x"73842b86",
   155 => x"a0712583",
   156 => x"7131700b",
   157 => x"0b0bbf80",
   158 => x"0c81712b",
   159 => x"ff05f688",
   160 => x"0cfdfc13",
   161 => x"ff122c78",
   162 => x"8829ff94",
   163 => x"0570812c",
   164 => x"80c39408",
   165 => x"52585255",
   166 => x"51525476",
   167 => x"802e8538",
   168 => x"70810751",
   169 => x"70f6940c",
   170 => x"71098105",
   171 => x"f6800c72",
   172 => x"098105f6",
   173 => x"840c0294",
   174 => x"050d0402",
   175 => x"f4050d74",
   176 => x"53727081",
   177 => x"055480f5",
   178 => x"2d527180",
   179 => x"2e893871",
   180 => x"5183842d",
   181 => x"85c10481",
   182 => x"0b80c2fc",
   183 => x"0c028c05",
   184 => x"0d0402f4",
   185 => x"050d7453",
   186 => x"80527173",
   187 => x"25913881",
   188 => x"808051c0",
   189 => x"115170fb",
   190 => x"38811252",
   191 => x"85ea0402",
   192 => x"8c050d04",
   193 => x"02f8050d",
   194 => x"e0528772",
   195 => x"0c84d851",
   196 => x"85e22d86",
   197 => x"720c0288",
   198 => x"050d0402",
   199 => x"fc050d80",
   200 => x"0bbf9c0c",
   201 => x"7251bac4",
   202 => x"2d028405",
   203 => x"0d0402fc",
   204 => x"050d810b",
   205 => x"bf9c0c72",
   206 => x"51bac42d",
   207 => x"0284050d",
   208 => x"0402ec05",
   209 => x"0d765580",
   210 => x"0bbf9c08",
   211 => x"54547281",
   212 => x"2e098106",
   213 => x"b6387452",
   214 => x"80c39851",
   215 => x"b1b22d80",
   216 => x"c2fc0874",
   217 => x"2ea53872",
   218 => x"73f40c54",
   219 => x"8a5185e2",
   220 => x"2d800bf4",
   221 => x"0c72bf98",
   222 => x"0c80c39c",
   223 => x"08bf940c",
   224 => x"800bbf90",
   225 => x"0c84800b",
   226 => x"bf8c0cbf",
   227 => x"9c08b238",
   228 => x"745280c3",
   229 => x"a451b1b2",
   230 => x"2d80c2fc",
   231 => x"08802ea1",
   232 => x"388170bf",
   233 => x"880c54ff",
   234 => x"0bbf840c",
   235 => x"80c3ac08",
   236 => x"80c3b40c",
   237 => x"80c1b808",
   238 => x"840780c1",
   239 => x"b80c87c6",
   240 => x"0473802e",
   241 => x"8d38bfa0",
   242 => x"5193d02d",
   243 => x"91c62d87",
   244 => x"d90480c0",
   245 => x"cc5193d0",
   246 => x"2d7380c2",
   247 => x"fc0c0294",
   248 => x"050d0402",
   249 => x"e4050d80",
   250 => x"70bf980c",
   251 => x"bf880c86",
   252 => x"0be00c90",
   253 => x"f72d8dc2",
   254 => x"2d81f92d",
   255 => x"83538151",
   256 => x"84a82dff",
   257 => x"13537280",
   258 => x"25f438bd",
   259 => x"b45185bb",
   260 => x"2da7f22d",
   261 => x"80c2fc08",
   262 => x"802e858f",
   263 => x"3886c151",
   264 => x"bae82dbf",
   265 => x"a05193d0",
   266 => x"2d91b22d",
   267 => x"8dce2d93",
   268 => x"e32d800b",
   269 => x"80c1b808",
   270 => x"70810655",
   271 => x"56567276",
   272 => x"2e833881",
   273 => x"56bfc00b",
   274 => x"80f52d70",
   275 => x"108e0677",
   276 => x"0776812a",
   277 => x"70810651",
   278 => x"55575472",
   279 => x"802e8538",
   280 => x"75900756",
   281 => x"bfd80b80",
   282 => x"f52d7085",
   283 => x"2ba00680",
   284 => x"c0880b80",
   285 => x"f52d7086",
   286 => x"2b81c006",
   287 => x"79730707",
   288 => x"78822a70",
   289 => x"81065157",
   290 => x"59525557",
   291 => x"72802e86",
   292 => x"38758280",
   293 => x"075675e4",
   294 => x"0c865380",
   295 => x"c2fc0883",
   296 => x"38845372",
   297 => x"e00cbf98",
   298 => x"08802e81",
   299 => x"8138bf8c",
   300 => x"0884802e",
   301 => x"09810680",
   302 => x"f53880c4",
   303 => x"845280c3",
   304 => x"9851b3ff",
   305 => x"2d80c2fc",
   306 => x"08802e91",
   307 => x"3880c484",
   308 => x"0b80c3b0",
   309 => x"0c800bbf",
   310 => x"8c0c89f2",
   311 => x"0486fada",
   312 => x"800bf80c",
   313 => x"86fada80",
   314 => x"0bfc0c80",
   315 => x"c2fc08bf",
   316 => x"980c80c3",
   317 => x"98085473",
   318 => x"b53880c4",
   319 => x"900b80f5",
   320 => x"2d537281",
   321 => x"2e098106",
   322 => x"a238820b",
   323 => x"f40c8aae",
   324 => x"04800bbf",
   325 => x"980c8b84",
   326 => x"0480c398",
   327 => x"51b3cf2d",
   328 => x"8b840480",
   329 => x"0bbf880c",
   330 => x"8c930473",
   331 => x"f40cbf98",
   332 => x"08802e80",
   333 => x"cf38ec08",
   334 => x"70810651",
   335 => x"5372802e",
   336 => x"80c23880",
   337 => x"c3b00884",
   338 => x"1180c3b0",
   339 => x"0c7008f0",
   340 => x"0c53bf94",
   341 => x"08fc0570",
   342 => x"bf940cbf",
   343 => x"90088405",
   344 => x"70bf900c",
   345 => x"71f80cfc",
   346 => x"0c538073",
   347 => x"25ffa238",
   348 => x"bf8c0884",
   349 => x"0570bf8c",
   350 => x"0c537284",
   351 => x"802eff99",
   352 => x"388ab604",
   353 => x"bf880880",
   354 => x"2efda138",
   355 => x"e408709f",
   356 => x"ff0671a0",
   357 => x"80065257",
   358 => x"5372802e",
   359 => x"80f93881",
   360 => x"0bec0c80",
   361 => x"e45185e2",
   362 => x"2d80c3b4",
   363 => x"0880c3ac",
   364 => x"0c800b80",
   365 => x"c3a40cbf",
   366 => x"8408802e",
   367 => x"953880c3",
   368 => x"a451b3cf",
   369 => x"2d80c3a4",
   370 => x"08bf8408",
   371 => x"2e098106",
   372 => x"ed38bf84",
   373 => x"088b0553",
   374 => x"80c3a408",
   375 => x"732eb438",
   376 => x"80c48455",
   377 => x"83fc54e8",
   378 => x"08757084",
   379 => x"05570cfc",
   380 => x"14547380",
   381 => x"25f13880",
   382 => x"c4845280",
   383 => x"c3a451b4",
   384 => x"a82d80c2",
   385 => x"fc08fe9b",
   386 => x"3880c3a4",
   387 => x"51b3cf2d",
   388 => x"8bd20480",
   389 => x"0bec0cbf",
   390 => x"8408762e",
   391 => x"fc8e3881",
   392 => x"0bec0c80",
   393 => x"e45185e2",
   394 => x"2d80c3b4",
   395 => x"0880c3ac",
   396 => x"0c800b80",
   397 => x"c3a40c75",
   398 => x"bf840c75",
   399 => x"802e9538",
   400 => x"80c3a451",
   401 => x"b3cf2d80",
   402 => x"c3a408bf",
   403 => x"84082e09",
   404 => x"8106ed38",
   405 => x"bf84088b",
   406 => x"055380c3",
   407 => x"a408732e",
   408 => x"80c23880",
   409 => x"c4845280",
   410 => x"c3a451b3",
   411 => x"ff2d80c2",
   412 => x"fc08802e",
   413 => x"9b3880c4",
   414 => x"845583fc",
   415 => x"54747084",
   416 => x"055608e8",
   417 => x"0cfc1454",
   418 => x"738025f1",
   419 => x"388d9a04",
   420 => x"80c2fc08",
   421 => x"bf880c8d",
   422 => x"a40480c3",
   423 => x"a451b3cf",
   424 => x"2d8cd404",
   425 => x"800bec0c",
   426 => x"88ac0480",
   427 => x"0b80c2fc",
   428 => x"0c029c05",
   429 => x"0d047198",
   430 => x"0c04ffb0",
   431 => x"0880c2fc",
   432 => x"0c04810b",
   433 => x"ffb00c04",
   434 => x"800bffb0",
   435 => x"0c0402f4",
   436 => x"050d80c3",
   437 => x"b8518fe1",
   438 => x"2dff0b80",
   439 => x"c2fc0825",
   440 => x"81883880",
   441 => x"c2fc0881",
   442 => x"f02e0981",
   443 => x"068a3881",
   444 => x"0b80c1b0",
   445 => x"0c8eea04",
   446 => x"80c2fc08",
   447 => x"81e02e09",
   448 => x"81068a38",
   449 => x"810b80c1",
   450 => x"b40c8eea",
   451 => x"0480c2fc",
   452 => x"085280c1",
   453 => x"b408802e",
   454 => x"893880c2",
   455 => x"fc088180",
   456 => x"05527184",
   457 => x"2c728f06",
   458 => x"535380c1",
   459 => x"b008802e",
   460 => x"9a387284",
   461 => x"2980c0f0",
   462 => x"05721381",
   463 => x"712b7009",
   464 => x"73080673",
   465 => x"0c515353",
   466 => x"8ede0472",
   467 => x"842980c0",
   468 => x"f0057213",
   469 => x"83712b72",
   470 => x"0807720c",
   471 => x"5353800b",
   472 => x"80c1b40c",
   473 => x"800b80c1",
   474 => x"b00c800b",
   475 => x"80c2fc0c",
   476 => x"028c050d",
   477 => x"0402f805",
   478 => x"0d80c0f0",
   479 => x"528f5180",
   480 => x"72708405",
   481 => x"540cff11",
   482 => x"51708025",
   483 => x"f2380288",
   484 => x"050d0402",
   485 => x"f0050d75",
   486 => x"518dc82d",
   487 => x"70822cfc",
   488 => x"0680c0f0",
   489 => x"1172109e",
   490 => x"06710870",
   491 => x"722a7083",
   492 => x"0682742b",
   493 => x"70097406",
   494 => x"760c5451",
   495 => x"56575351",
   496 => x"538dc22d",
   497 => x"7180c2fc",
   498 => x"0c029005",
   499 => x"0d0402fc",
   500 => x"050d7251",
   501 => x"80710c80",
   502 => x"0b84120c",
   503 => x"0284050d",
   504 => x"0402f005",
   505 => x"0d757008",
   506 => x"84120853",
   507 => x"5353ff54",
   508 => x"71712ea8",
   509 => x"388dc82d",
   510 => x"84130870",
   511 => x"84291488",
   512 => x"11700870",
   513 => x"81ff0684",
   514 => x"18088111",
   515 => x"8706841a",
   516 => x"0c535155",
   517 => x"5151518d",
   518 => x"c22d7154",
   519 => x"7380c2fc",
   520 => x"0c029005",
   521 => x"0d0402f4",
   522 => x"050d8dc8",
   523 => x"2de00870",
   524 => x"8b2a7081",
   525 => x"06515253",
   526 => x"70802ea1",
   527 => x"3880c3b8",
   528 => x"08708429",
   529 => x"80c3c005",
   530 => x"7481ff06",
   531 => x"710c5151",
   532 => x"80c3b808",
   533 => x"81118706",
   534 => x"80c3b80c",
   535 => x"51728c2c",
   536 => x"bf0680c3",
   537 => x"e00c800b",
   538 => x"80c3e40c",
   539 => x"8dba2d8d",
   540 => x"c22d028c",
   541 => x"050d0402",
   542 => x"fc050d80",
   543 => x"c3b8518f",
   544 => x"ce2d8ef5",
   545 => x"2d90a651",
   546 => x"8db62d02",
   547 => x"84050d04",
   548 => x"02f8050d",
   549 => x"8fcf5281",
   550 => x"5185e22d",
   551 => x"ff125271",
   552 => x"8025f438",
   553 => x"0288050d",
   554 => x"0480c3f0",
   555 => x"0880c2fc",
   556 => x"0c0402fc",
   557 => x"050d810b",
   558 => x"80c1bc0c",
   559 => x"815184a8",
   560 => x"2d028405",
   561 => x"0d0402fc",
   562 => x"050d91d0",
   563 => x"048dce2d",
   564 => x"80f6518f",
   565 => x"932d80c2",
   566 => x"fc08f238",
   567 => x"80da518f",
   568 => x"932d80c2",
   569 => x"fc08e638",
   570 => x"80c2fc08",
   571 => x"80c1bc0c",
   572 => x"80c2fc08",
   573 => x"5184a82d",
   574 => x"0284050d",
   575 => x"0402ec05",
   576 => x"0d765480",
   577 => x"52870b88",
   578 => x"1580f52d",
   579 => x"56537472",
   580 => x"248338a0",
   581 => x"53725183",
   582 => x"842d8112",
   583 => x"8b1580f5",
   584 => x"2d545272",
   585 => x"7225de38",
   586 => x"0294050d",
   587 => x"0402f005",
   588 => x"0d80c3f0",
   589 => x"085481f9",
   590 => x"2d800b80",
   591 => x"c3f40c73",
   592 => x"08802e81",
   593 => x"8638820b",
   594 => x"80c3900c",
   595 => x"80c3f408",
   596 => x"8f0680c3",
   597 => x"8c0c7308",
   598 => x"5271832e",
   599 => x"96387183",
   600 => x"26893871",
   601 => x"812eaf38",
   602 => x"93b40471",
   603 => x"852e9f38",
   604 => x"93b40488",
   605 => x"1480f52d",
   606 => x"841508bd",
   607 => x"cc535452",
   608 => x"85bb2d71",
   609 => x"84291370",
   610 => x"08525293",
   611 => x"b8047351",
   612 => x"91fd2d93",
   613 => x"b40480c1",
   614 => x"b8088815",
   615 => x"082c7081",
   616 => x"06515271",
   617 => x"802e8738",
   618 => x"bdd05193",
   619 => x"b104bdd4",
   620 => x"5185bb2d",
   621 => x"84140851",
   622 => x"85bb2d80",
   623 => x"c3f40881",
   624 => x"0580c3f4",
   625 => x"0c8c1454",
   626 => x"92bf0402",
   627 => x"90050d04",
   628 => x"7180c3f0",
   629 => x"0c92ad2d",
   630 => x"80c3f408",
   631 => x"ff0580c3",
   632 => x"f80c0402",
   633 => x"e8050d80",
   634 => x"c3f00880",
   635 => x"c3fc0857",
   636 => x"5580f651",
   637 => x"8f932d80",
   638 => x"c2fc0881",
   639 => x"2a708106",
   640 => x"51527180",
   641 => x"2ea23894",
   642 => x"8d048dce",
   643 => x"2d80f651",
   644 => x"8f932d80",
   645 => x"c2fc08f2",
   646 => x"3880c1bc",
   647 => x"08813270",
   648 => x"80c1bc0c",
   649 => x"5184a82d",
   650 => x"80c3e008",
   651 => x"a0065280",
   652 => x"72259838",
   653 => x"91902d8d",
   654 => x"ce2d80c1",
   655 => x"bc088132",
   656 => x"7080c1bc",
   657 => x"0c705252",
   658 => x"84a82d80",
   659 => x"0b80c3e8",
   660 => x"0c800b80",
   661 => x"c3ec0c80",
   662 => x"c1bc0883",
   663 => x"8d3880da",
   664 => x"518f932d",
   665 => x"80c2fc08",
   666 => x"802e8c38",
   667 => x"80c3e808",
   668 => x"81800780",
   669 => x"c3e80c80",
   670 => x"d9518f93",
   671 => x"2d80c2fc",
   672 => x"08802e8c",
   673 => x"3880c3e8",
   674 => x"0880c007",
   675 => x"80c3e80c",
   676 => x"8194518f",
   677 => x"932d80c2",
   678 => x"fc08802e",
   679 => x"8b3880c3",
   680 => x"e8089007",
   681 => x"80c3e80c",
   682 => x"8191518f",
   683 => x"932d80c2",
   684 => x"fc08802e",
   685 => x"8b3880c3",
   686 => x"e808a007",
   687 => x"80c3e80c",
   688 => x"81f5518f",
   689 => x"932d80c2",
   690 => x"fc08802e",
   691 => x"8b3880c3",
   692 => x"e8088107",
   693 => x"80c3e80c",
   694 => x"81f2518f",
   695 => x"932d80c2",
   696 => x"fc08802e",
   697 => x"8b3880c3",
   698 => x"e8088207",
   699 => x"80c3e80c",
   700 => x"81eb518f",
   701 => x"932d80c2",
   702 => x"fc08802e",
   703 => x"8b3880c3",
   704 => x"e8088407",
   705 => x"80c3e80c",
   706 => x"81f4518f",
   707 => x"932d80c2",
   708 => x"fc08802e",
   709 => x"8b3880c3",
   710 => x"e8088807",
   711 => x"80c3e80c",
   712 => x"80d8518f",
   713 => x"932d80c2",
   714 => x"fc08802e",
   715 => x"8c3880c3",
   716 => x"ec088180",
   717 => x"0780c3ec",
   718 => x"0c92518f",
   719 => x"932d80c2",
   720 => x"fc08802e",
   721 => x"8c3880c3",
   722 => x"ec0880c0",
   723 => x"0780c3ec",
   724 => x"0c94518f",
   725 => x"932d80c2",
   726 => x"fc08802e",
   727 => x"8b3880c3",
   728 => x"ec089007",
   729 => x"80c3ec0c",
   730 => x"91518f93",
   731 => x"2d80c2fc",
   732 => x"08802e8b",
   733 => x"3880c3ec",
   734 => x"08a00780",
   735 => x"c3ec0c9d",
   736 => x"518f932d",
   737 => x"80c2fc08",
   738 => x"802e8b38",
   739 => x"80c3ec08",
   740 => x"810780c3",
   741 => x"ec0c9b51",
   742 => x"8f932d80",
   743 => x"c2fc0880",
   744 => x"2e8b3880",
   745 => x"c3ec0882",
   746 => x"0780c3ec",
   747 => x"0c9c518f",
   748 => x"932d80c2",
   749 => x"fc08802e",
   750 => x"8b3880c3",
   751 => x"ec088407",
   752 => x"80c3ec0c",
   753 => x"a3518f93",
   754 => x"2d80c2fc",
   755 => x"08802e8b",
   756 => x"3880c3ec",
   757 => x"08880780",
   758 => x"c3ec0c81",
   759 => x"fd518f93",
   760 => x"2d81fa51",
   761 => x"8f932d9e",
   762 => x"8c0481f5",
   763 => x"518f932d",
   764 => x"80c2fc08",
   765 => x"812a7081",
   766 => x"06515271",
   767 => x"8e3880c3",
   768 => x"e0089006",
   769 => x"52807225",
   770 => x"80c23880",
   771 => x"c3e00890",
   772 => x"06528072",
   773 => x"25843891",
   774 => x"902d80c3",
   775 => x"f8085271",
   776 => x"802e8a38",
   777 => x"ff1280c3",
   778 => x"f80c98cc",
   779 => x"0480c3f4",
   780 => x"081080c3",
   781 => x"f4080570",
   782 => x"84291651",
   783 => x"52881208",
   784 => x"802e8938",
   785 => x"ff518812",
   786 => x"0852712d",
   787 => x"81f2518f",
   788 => x"932d80c2",
   789 => x"fc08812a",
   790 => x"70810651",
   791 => x"52718e38",
   792 => x"80c3e008",
   793 => x"88065280",
   794 => x"722580c3",
   795 => x"3880c3e0",
   796 => x"08880652",
   797 => x"80722584",
   798 => x"3891902d",
   799 => x"80c3f408",
   800 => x"ff1180c3",
   801 => x"f8085653",
   802 => x"53737225",
   803 => x"8a388114",
   804 => x"80c3f80c",
   805 => x"99af0472",
   806 => x"10137084",
   807 => x"29165152",
   808 => x"88120880",
   809 => x"2e8938fe",
   810 => x"51881208",
   811 => x"52712d81",
   812 => x"fd518f93",
   813 => x"2d80c2fc",
   814 => x"08812a70",
   815 => x"81065152",
   816 => x"71802eb1",
   817 => x"3880c3f8",
   818 => x"08802e8a",
   819 => x"38800b80",
   820 => x"c3f80c99",
   821 => x"f50480c3",
   822 => x"f4081080",
   823 => x"c3f40805",
   824 => x"70842916",
   825 => x"51528812",
   826 => x"08802e89",
   827 => x"38fd5188",
   828 => x"12085271",
   829 => x"2d81fa51",
   830 => x"8f932d80",
   831 => x"c2fc0881",
   832 => x"2a708106",
   833 => x"51527180",
   834 => x"2eb13880",
   835 => x"c3f408ff",
   836 => x"11545280",
   837 => x"c3f80873",
   838 => x"25893872",
   839 => x"80c3f80c",
   840 => x"9abb0471",
   841 => x"10127084",
   842 => x"29165152",
   843 => x"88120880",
   844 => x"2e8938fc",
   845 => x"51881208",
   846 => x"52712d80",
   847 => x"c3f80870",
   848 => x"53547380",
   849 => x"2e8a388c",
   850 => x"15ff1555",
   851 => x"559ac204",
   852 => x"820b80c3",
   853 => x"900c718f",
   854 => x"0680c38c",
   855 => x"0c81eb51",
   856 => x"8f932d80",
   857 => x"c2fc0881",
   858 => x"2a708106",
   859 => x"51527180",
   860 => x"2ead3874",
   861 => x"08852e09",
   862 => x"8106a438",
   863 => x"881580f5",
   864 => x"2dff0552",
   865 => x"71881681",
   866 => x"b72d7198",
   867 => x"2b527180",
   868 => x"25883880",
   869 => x"0b881681",
   870 => x"b72d7451",
   871 => x"91fd2d81",
   872 => x"f4518f93",
   873 => x"2d80c2fc",
   874 => x"08812a70",
   875 => x"81065152",
   876 => x"71802eb3",
   877 => x"38740885",
   878 => x"2e098106",
   879 => x"aa388815",
   880 => x"80f52d81",
   881 => x"05527188",
   882 => x"1681b72d",
   883 => x"7181ff06",
   884 => x"8b1680f5",
   885 => x"2d545272",
   886 => x"72278738",
   887 => x"72881681",
   888 => x"b72d7451",
   889 => x"91fd2d80",
   890 => x"da518f93",
   891 => x"2d80c2fc",
   892 => x"08812a70",
   893 => x"81065152",
   894 => x"718e3880",
   895 => x"c3e00881",
   896 => x"06528072",
   897 => x"2581bc38",
   898 => x"80c3f008",
   899 => x"80c3e008",
   900 => x"81065353",
   901 => x"80722584",
   902 => x"3891902d",
   903 => x"80c3f808",
   904 => x"5473802e",
   905 => x"8a388c13",
   906 => x"ff155553",
   907 => x"9ca10472",
   908 => x"08527182",
   909 => x"2ea63871",
   910 => x"82268938",
   911 => x"71812eaa",
   912 => x"389dc304",
   913 => x"71832eb4",
   914 => x"3871842e",
   915 => x"09810680",
   916 => x"f2388813",
   917 => x"085193d0",
   918 => x"2d9dc304",
   919 => x"80c3f808",
   920 => x"51881308",
   921 => x"52712d9d",
   922 => x"c304810b",
   923 => x"8814082b",
   924 => x"80c1b808",
   925 => x"3280c1b8",
   926 => x"0c9d9704",
   927 => x"881380f5",
   928 => x"2d81058b",
   929 => x"1480f52d",
   930 => x"53547174",
   931 => x"24833880",
   932 => x"54738814",
   933 => x"81b72d92",
   934 => x"ad2d9dc3",
   935 => x"04750880",
   936 => x"2ea43875",
   937 => x"08518f93",
   938 => x"2d80c2fc",
   939 => x"08810652",
   940 => x"71802e8c",
   941 => x"3880c3f8",
   942 => x"08518416",
   943 => x"0852712d",
   944 => x"88165675",
   945 => x"d8388054",
   946 => x"800b80c3",
   947 => x"900c738f",
   948 => x"0680c38c",
   949 => x"0ca05273",
   950 => x"80c3f808",
   951 => x"2e098106",
   952 => x"993880c3",
   953 => x"f408ff05",
   954 => x"74327009",
   955 => x"81057072",
   956 => x"079f2a91",
   957 => x"71315151",
   958 => x"53537151",
   959 => x"83842d81",
   960 => x"14548e74",
   961 => x"25c23880",
   962 => x"c1bc0852",
   963 => x"7180c2fc",
   964 => x"0c029805",
   965 => x"0d0402f4",
   966 => x"050dd452",
   967 => x"81ff720c",
   968 => x"71085381",
   969 => x"ff720c72",
   970 => x"882b83fe",
   971 => x"80067208",
   972 => x"7081ff06",
   973 => x"51525381",
   974 => x"ff720c72",
   975 => x"7107882b",
   976 => x"72087081",
   977 => x"ff065152",
   978 => x"5381ff72",
   979 => x"0c727107",
   980 => x"882b7208",
   981 => x"7081ff06",
   982 => x"720780c2",
   983 => x"fc0c5253",
   984 => x"028c050d",
   985 => x"0402f405",
   986 => x"0d747671",
   987 => x"81ff06d4",
   988 => x"0c535380",
   989 => x"c4800885",
   990 => x"3871892b",
   991 => x"5271982a",
   992 => x"d40c7190",
   993 => x"2a7081ff",
   994 => x"06d40c51",
   995 => x"71882a70",
   996 => x"81ff06d4",
   997 => x"0c517181",
   998 => x"ff06d40c",
   999 => x"72902a70",
  1000 => x"81ff06d4",
  1001 => x"0c51d408",
  1002 => x"7081ff06",
  1003 => x"515182b8",
  1004 => x"bf527081",
  1005 => x"ff2e0981",
  1006 => x"06943881",
  1007 => x"ff0bd40c",
  1008 => x"d4087081",
  1009 => x"ff06ff14",
  1010 => x"54515171",
  1011 => x"e5387080",
  1012 => x"c2fc0c02",
  1013 => x"8c050d04",
  1014 => x"02fc050d",
  1015 => x"81c75181",
  1016 => x"ff0bd40c",
  1017 => x"ff115170",
  1018 => x"8025f438",
  1019 => x"0284050d",
  1020 => x"0402f405",
  1021 => x"0d81ff0b",
  1022 => x"d40c9353",
  1023 => x"805287fc",
  1024 => x"80c1519e",
  1025 => x"e52d80c2",
  1026 => x"fc088b38",
  1027 => x"81ff0bd4",
  1028 => x"0c8153a0",
  1029 => x"9f049fd8",
  1030 => x"2dff1353",
  1031 => x"72de3872",
  1032 => x"80c2fc0c",
  1033 => x"028c050d",
  1034 => x"0402ec05",
  1035 => x"0d810b80",
  1036 => x"c4800c84",
  1037 => x"54d00870",
  1038 => x"8f2a7081",
  1039 => x"06515153",
  1040 => x"72f33872",
  1041 => x"d00c9fd8",
  1042 => x"2dbdd851",
  1043 => x"85bb2dd0",
  1044 => x"08708f2a",
  1045 => x"70810651",
  1046 => x"515372f3",
  1047 => x"38810bd0",
  1048 => x"0cb15380",
  1049 => x"5284d480",
  1050 => x"c0519ee5",
  1051 => x"2d80c2fc",
  1052 => x"08812e93",
  1053 => x"3872822e",
  1054 => x"bf38ff13",
  1055 => x"5372e438",
  1056 => x"ff145473",
  1057 => x"ffaf389f",
  1058 => x"d82d83aa",
  1059 => x"52849c80",
  1060 => x"c8519ee5",
  1061 => x"2d80c2fc",
  1062 => x"08812e09",
  1063 => x"81069338",
  1064 => x"9e962d80",
  1065 => x"c2fc0883",
  1066 => x"ffff0653",
  1067 => x"7283aa2e",
  1068 => x"9d389ff1",
  1069 => x"2da1c904",
  1070 => x"bde45185",
  1071 => x"bb2d8053",
  1072 => x"a39e04bd",
  1073 => x"fc5185bb",
  1074 => x"2d8054a2",
  1075 => x"ef0481ff",
  1076 => x"0bd40cb1",
  1077 => x"549fd82d",
  1078 => x"8fcf5380",
  1079 => x"5287fc80",
  1080 => x"f7519ee5",
  1081 => x"2d80c2fc",
  1082 => x"085580c2",
  1083 => x"fc08812e",
  1084 => x"0981069c",
  1085 => x"3881ff0b",
  1086 => x"d40c820a",
  1087 => x"52849c80",
  1088 => x"e9519ee5",
  1089 => x"2d80c2fc",
  1090 => x"08802e8d",
  1091 => x"389fd82d",
  1092 => x"ff135372",
  1093 => x"c638a2e2",
  1094 => x"0481ff0b",
  1095 => x"d40c80c2",
  1096 => x"fc085287",
  1097 => x"fc80fa51",
  1098 => x"9ee52d80",
  1099 => x"c2fc08b2",
  1100 => x"3881ff0b",
  1101 => x"d40cd408",
  1102 => x"5381ff0b",
  1103 => x"d40c81ff",
  1104 => x"0bd40c81",
  1105 => x"ff0bd40c",
  1106 => x"81ff0bd4",
  1107 => x"0c72862a",
  1108 => x"70810676",
  1109 => x"56515372",
  1110 => x"963880c2",
  1111 => x"fc0854a2",
  1112 => x"ef047382",
  1113 => x"2efedc38",
  1114 => x"ff145473",
  1115 => x"fee73873",
  1116 => x"80c4800c",
  1117 => x"738b3881",
  1118 => x"5287fc80",
  1119 => x"d0519ee5",
  1120 => x"2d81ff0b",
  1121 => x"d40cd008",
  1122 => x"708f2a70",
  1123 => x"81065151",
  1124 => x"5372f338",
  1125 => x"72d00c81",
  1126 => x"ff0bd40c",
  1127 => x"81537280",
  1128 => x"c2fc0c02",
  1129 => x"94050d04",
  1130 => x"02e8050d",
  1131 => x"785681ff",
  1132 => x"0bd40cd0",
  1133 => x"08708f2a",
  1134 => x"70810651",
  1135 => x"515372f3",
  1136 => x"3882810b",
  1137 => x"d00c81ff",
  1138 => x"0bd40c77",
  1139 => x"5287fc80",
  1140 => x"d8519ee5",
  1141 => x"2d80c2fc",
  1142 => x"08802e8c",
  1143 => x"38be8c51",
  1144 => x"85bb2d81",
  1145 => x"53a4e004",
  1146 => x"81ff0bd4",
  1147 => x"0c81fe0b",
  1148 => x"d40c80ff",
  1149 => x"55757084",
  1150 => x"05570870",
  1151 => x"982ad40c",
  1152 => x"70902c70",
  1153 => x"81ff06d4",
  1154 => x"0c547088",
  1155 => x"2c7081ff",
  1156 => x"06d40c54",
  1157 => x"7081ff06",
  1158 => x"d40c54ff",
  1159 => x"15557480",
  1160 => x"25d33881",
  1161 => x"ff0bd40c",
  1162 => x"81ff0bd4",
  1163 => x"0c81ff0b",
  1164 => x"d40c868d",
  1165 => x"a05481ff",
  1166 => x"0bd40cd4",
  1167 => x"0881ff06",
  1168 => x"55748738",
  1169 => x"ff145473",
  1170 => x"ed3881ff",
  1171 => x"0bd40cd0",
  1172 => x"08708f2a",
  1173 => x"70810651",
  1174 => x"515372f3",
  1175 => x"3872d00c",
  1176 => x"7280c2fc",
  1177 => x"0c029805",
  1178 => x"0d0402e8",
  1179 => x"050d7855",
  1180 => x"805681ff",
  1181 => x"0bd40cd0",
  1182 => x"08708f2a",
  1183 => x"70810651",
  1184 => x"515372f3",
  1185 => x"3882810b",
  1186 => x"d00c81ff",
  1187 => x"0bd40c77",
  1188 => x"5287fc80",
  1189 => x"d1519ee5",
  1190 => x"2d80dbc6",
  1191 => x"df5480c2",
  1192 => x"fc08802e",
  1193 => x"8a38be9c",
  1194 => x"5185bb2d",
  1195 => x"a6830481",
  1196 => x"ff0bd40c",
  1197 => x"d4087081",
  1198 => x"ff065153",
  1199 => x"7281fe2e",
  1200 => x"0981069e",
  1201 => x"3880ff53",
  1202 => x"9e962d80",
  1203 => x"c2fc0875",
  1204 => x"70840557",
  1205 => x"0cff1353",
  1206 => x"728025ec",
  1207 => x"388156a5",
  1208 => x"e804ff14",
  1209 => x"5473c838",
  1210 => x"81ff0bd4",
  1211 => x"0c81ff0b",
  1212 => x"d40cd008",
  1213 => x"708f2a70",
  1214 => x"81065151",
  1215 => x"5372f338",
  1216 => x"72d00c75",
  1217 => x"80c2fc0c",
  1218 => x"0298050d",
  1219 => x"0402e805",
  1220 => x"0d77797b",
  1221 => x"58555580",
  1222 => x"53727625",
  1223 => x"a3387470",
  1224 => x"81055680",
  1225 => x"f52d7470",
  1226 => x"81055680",
  1227 => x"f52d5252",
  1228 => x"71712e86",
  1229 => x"388151a6",
  1230 => x"c2048113",
  1231 => x"53a69904",
  1232 => x"80517080",
  1233 => x"c2fc0c02",
  1234 => x"98050d04",
  1235 => x"02ec050d",
  1236 => x"76557480",
  1237 => x"2e80c238",
  1238 => x"9a1580e0",
  1239 => x"2d51b582",
  1240 => x"2d80c2fc",
  1241 => x"0880c2fc",
  1242 => x"0880cab4",
  1243 => x"0c80c2fc",
  1244 => x"08545480",
  1245 => x"ca900880",
  1246 => x"2e9a3894",
  1247 => x"1580e02d",
  1248 => x"51b5822d",
  1249 => x"80c2fc08",
  1250 => x"902b83ff",
  1251 => x"f00a0670",
  1252 => x"75075153",
  1253 => x"7280cab4",
  1254 => x"0c80cab4",
  1255 => x"08537280",
  1256 => x"2e9d3880",
  1257 => x"ca8808fe",
  1258 => x"14712980",
  1259 => x"ca9c0805",
  1260 => x"80cab80c",
  1261 => x"70842b80",
  1262 => x"ca940c54",
  1263 => x"a7ed0480",
  1264 => x"caa00880",
  1265 => x"cab40c80",
  1266 => x"caa40880",
  1267 => x"cab80c80",
  1268 => x"ca900880",
  1269 => x"2e8b3880",
  1270 => x"ca880884",
  1271 => x"2b53a7e8",
  1272 => x"0480caa8",
  1273 => x"08842b53",
  1274 => x"7280ca94",
  1275 => x"0c029405",
  1276 => x"0d0402d8",
  1277 => x"050d800b",
  1278 => x"80ca900c",
  1279 => x"8454a0a9",
  1280 => x"2d80c2fc",
  1281 => x"08802e97",
  1282 => x"3880c484",
  1283 => x"528051a4",
  1284 => x"ea2d80c2",
  1285 => x"fc08802e",
  1286 => x"8638fe54",
  1287 => x"a8a704ff",
  1288 => x"14547380",
  1289 => x"24d83873",
  1290 => x"8c38beac",
  1291 => x"5185bb2d",
  1292 => x"7355adf4",
  1293 => x"04805681",
  1294 => x"0b80cabc",
  1295 => x"0c8853be",
  1296 => x"c05280c4",
  1297 => x"ba51a68d",
  1298 => x"2d80c2fc",
  1299 => x"08762e09",
  1300 => x"81068938",
  1301 => x"80c2fc08",
  1302 => x"80cabc0c",
  1303 => x"8853becc",
  1304 => x"5280c4d6",
  1305 => x"51a68d2d",
  1306 => x"80c2fc08",
  1307 => x"893880c2",
  1308 => x"fc0880ca",
  1309 => x"bc0c80ca",
  1310 => x"bc08802e",
  1311 => x"81803880",
  1312 => x"c7ca0b80",
  1313 => x"f52d80c7",
  1314 => x"cb0b80f5",
  1315 => x"2d71982b",
  1316 => x"71902b07",
  1317 => x"80c7cc0b",
  1318 => x"80f52d70",
  1319 => x"882b7207",
  1320 => x"80c7cd0b",
  1321 => x"80f52d71",
  1322 => x"0780c882",
  1323 => x"0b80f52d",
  1324 => x"80c8830b",
  1325 => x"80f52d71",
  1326 => x"882b0753",
  1327 => x"5f54525a",
  1328 => x"56575573",
  1329 => x"81abaa2e",
  1330 => x"0981068e",
  1331 => x"387551b4",
  1332 => x"d12d80c2",
  1333 => x"fc0856a9",
  1334 => x"e7047382",
  1335 => x"d4d52e87",
  1336 => x"38bed851",
  1337 => x"aab00480",
  1338 => x"c4845275",
  1339 => x"51a4ea2d",
  1340 => x"80c2fc08",
  1341 => x"5580c2fc",
  1342 => x"08802e83",
  1343 => x"f7388853",
  1344 => x"becc5280",
  1345 => x"c4d651a6",
  1346 => x"8d2d80c2",
  1347 => x"fc088a38",
  1348 => x"810b80ca",
  1349 => x"900caab6",
  1350 => x"048853be",
  1351 => x"c05280c4",
  1352 => x"ba51a68d",
  1353 => x"2d80c2fc",
  1354 => x"08802e8a",
  1355 => x"38beec51",
  1356 => x"85bb2dab",
  1357 => x"950480c8",
  1358 => x"820b80f5",
  1359 => x"2d547380",
  1360 => x"d52e0981",
  1361 => x"0680ce38",
  1362 => x"80c8830b",
  1363 => x"80f52d54",
  1364 => x"7381aa2e",
  1365 => x"098106bd",
  1366 => x"38800b80",
  1367 => x"c4840b80",
  1368 => x"f52d5654",
  1369 => x"7481e92e",
  1370 => x"83388154",
  1371 => x"7481eb2e",
  1372 => x"8c388055",
  1373 => x"73752e09",
  1374 => x"810682f8",
  1375 => x"3880c48f",
  1376 => x"0b80f52d",
  1377 => x"55748e38",
  1378 => x"80c4900b",
  1379 => x"80f52d54",
  1380 => x"73822e86",
  1381 => x"388055ad",
  1382 => x"f40480c4",
  1383 => x"910b80f5",
  1384 => x"2d7080ca",
  1385 => x"880cff05",
  1386 => x"80ca8c0c",
  1387 => x"80c4920b",
  1388 => x"80f52d80",
  1389 => x"c4930b80",
  1390 => x"f52d5876",
  1391 => x"05778280",
  1392 => x"29057080",
  1393 => x"ca980c80",
  1394 => x"c4940b80",
  1395 => x"f52d7080",
  1396 => x"caac0c80",
  1397 => x"ca900859",
  1398 => x"57587680",
  1399 => x"2e81b638",
  1400 => x"8853becc",
  1401 => x"5280c4d6",
  1402 => x"51a68d2d",
  1403 => x"80c2fc08",
  1404 => x"82823880",
  1405 => x"ca880870",
  1406 => x"842b80ca",
  1407 => x"940c7080",
  1408 => x"caa80c80",
  1409 => x"c4a90b80",
  1410 => x"f52d80c4",
  1411 => x"a80b80f5",
  1412 => x"2d718280",
  1413 => x"290580c4",
  1414 => x"aa0b80f5",
  1415 => x"2d708480",
  1416 => x"80291280",
  1417 => x"c4ab0b80",
  1418 => x"f52d7081",
  1419 => x"800a2912",
  1420 => x"7080cab0",
  1421 => x"0c80caac",
  1422 => x"08712980",
  1423 => x"ca980805",
  1424 => x"7080ca9c",
  1425 => x"0c80c4b1",
  1426 => x"0b80f52d",
  1427 => x"80c4b00b",
  1428 => x"80f52d71",
  1429 => x"82802905",
  1430 => x"80c4b20b",
  1431 => x"80f52d70",
  1432 => x"84808029",
  1433 => x"1280c4b3",
  1434 => x"0b80f52d",
  1435 => x"70982b81",
  1436 => x"f00a0672",
  1437 => x"057080ca",
  1438 => x"a00cfe11",
  1439 => x"7e297705",
  1440 => x"80caa40c",
  1441 => x"52595243",
  1442 => x"545e5152",
  1443 => x"59525d57",
  1444 => x"5957aded",
  1445 => x"0480c496",
  1446 => x"0b80f52d",
  1447 => x"80c4950b",
  1448 => x"80f52d71",
  1449 => x"82802905",
  1450 => x"7080ca94",
  1451 => x"0c70a029",
  1452 => x"83ff0570",
  1453 => x"892a7080",
  1454 => x"caa80c80",
  1455 => x"c49b0b80",
  1456 => x"f52d80c4",
  1457 => x"9a0b80f5",
  1458 => x"2d718280",
  1459 => x"29057080",
  1460 => x"cab00c7b",
  1461 => x"71291e70",
  1462 => x"80caa40c",
  1463 => x"7d80caa0",
  1464 => x"0c730580",
  1465 => x"ca9c0c55",
  1466 => x"5e515155",
  1467 => x"558051a6",
  1468 => x"cc2d8155",
  1469 => x"7480c2fc",
  1470 => x"0c02a805",
  1471 => x"0d0402ec",
  1472 => x"050d7670",
  1473 => x"872c7180",
  1474 => x"ff065556",
  1475 => x"5480ca90",
  1476 => x"088a3873",
  1477 => x"882c7481",
  1478 => x"ff065455",
  1479 => x"80c48452",
  1480 => x"80ca9808",
  1481 => x"1551a4ea",
  1482 => x"2d80c2fc",
  1483 => x"085480c2",
  1484 => x"fc08802e",
  1485 => x"b83880ca",
  1486 => x"9008802e",
  1487 => x"9a387284",
  1488 => x"2980c484",
  1489 => x"05700852",
  1490 => x"53b4d12d",
  1491 => x"80c2fc08",
  1492 => x"f00a0653",
  1493 => x"aeeb0472",
  1494 => x"1080c484",
  1495 => x"057080e0",
  1496 => x"2d5253b5",
  1497 => x"822d80c2",
  1498 => x"fc085372",
  1499 => x"547380c2",
  1500 => x"fc0c0294",
  1501 => x"050d0402",
  1502 => x"e0050d79",
  1503 => x"70842c80",
  1504 => x"cab80805",
  1505 => x"718f0652",
  1506 => x"5553728a",
  1507 => x"3880c484",
  1508 => x"527351a4",
  1509 => x"ea2d72a0",
  1510 => x"2980c484",
  1511 => x"05548074",
  1512 => x"80f52d56",
  1513 => x"5374732e",
  1514 => x"83388153",
  1515 => x"7481e52e",
  1516 => x"81f43881",
  1517 => x"70740654",
  1518 => x"5872802e",
  1519 => x"81e8388b",
  1520 => x"1480f52d",
  1521 => x"70832a79",
  1522 => x"06585676",
  1523 => x"9b3880c1",
  1524 => x"c0085372",
  1525 => x"89387280",
  1526 => x"c8840b81",
  1527 => x"b72d7680",
  1528 => x"c1c00c73",
  1529 => x"53b1a804",
  1530 => x"758f2e09",
  1531 => x"810681b6",
  1532 => x"38749f06",
  1533 => x"8d2980c7",
  1534 => x"f7115153",
  1535 => x"811480f5",
  1536 => x"2d737081",
  1537 => x"055581b7",
  1538 => x"2d831480",
  1539 => x"f52d7370",
  1540 => x"81055581",
  1541 => x"b72d8514",
  1542 => x"80f52d73",
  1543 => x"70810555",
  1544 => x"81b72d87",
  1545 => x"1480f52d",
  1546 => x"73708105",
  1547 => x"5581b72d",
  1548 => x"891480f5",
  1549 => x"2d737081",
  1550 => x"055581b7",
  1551 => x"2d8e1480",
  1552 => x"f52d7370",
  1553 => x"81055581",
  1554 => x"b72d9014",
  1555 => x"80f52d73",
  1556 => x"70810555",
  1557 => x"81b72d92",
  1558 => x"1480f52d",
  1559 => x"73708105",
  1560 => x"5581b72d",
  1561 => x"941480f5",
  1562 => x"2d737081",
  1563 => x"055581b7",
  1564 => x"2d961480",
  1565 => x"f52d7370",
  1566 => x"81055581",
  1567 => x"b72d9814",
  1568 => x"80f52d73",
  1569 => x"70810555",
  1570 => x"81b72d9c",
  1571 => x"1480f52d",
  1572 => x"73708105",
  1573 => x"5581b72d",
  1574 => x"9e1480f5",
  1575 => x"2d7381b7",
  1576 => x"2d7780c1",
  1577 => x"c00c8053",
  1578 => x"7280c2fc",
  1579 => x"0c02a005",
  1580 => x"0d0402cc",
  1581 => x"050d7e60",
  1582 => x"5e5a800b",
  1583 => x"80cab408",
  1584 => x"80cab808",
  1585 => x"595c5680",
  1586 => x"5880ca94",
  1587 => x"08782e81",
  1588 => x"b838778f",
  1589 => x"06a01757",
  1590 => x"54739138",
  1591 => x"80c48452",
  1592 => x"76518117",
  1593 => x"57a4ea2d",
  1594 => x"80c48456",
  1595 => x"807680f5",
  1596 => x"2d565474",
  1597 => x"742e8338",
  1598 => x"81547481",
  1599 => x"e52e80fd",
  1600 => x"38817075",
  1601 => x"06555c73",
  1602 => x"802e80f1",
  1603 => x"388b1680",
  1604 => x"f52d9806",
  1605 => x"597880e5",
  1606 => x"388b537c",
  1607 => x"527551a6",
  1608 => x"8d2d80c2",
  1609 => x"fc0880d5",
  1610 => x"389c1608",
  1611 => x"51b4d12d",
  1612 => x"80c2fc08",
  1613 => x"841b0c9a",
  1614 => x"1680e02d",
  1615 => x"51b5822d",
  1616 => x"80c2fc08",
  1617 => x"80c2fc08",
  1618 => x"881c0c80",
  1619 => x"c2fc0855",
  1620 => x"5580ca90",
  1621 => x"08802e99",
  1622 => x"38941680",
  1623 => x"e02d51b5",
  1624 => x"822d80c2",
  1625 => x"fc08902b",
  1626 => x"83fff00a",
  1627 => x"06701651",
  1628 => x"5473881b",
  1629 => x"0c787a0c",
  1630 => x"7b54b3c5",
  1631 => x"04811858",
  1632 => x"80ca9408",
  1633 => x"7826feca",
  1634 => x"3880ca90",
  1635 => x"08802eb3",
  1636 => x"387a51ad",
  1637 => x"fe2d80c2",
  1638 => x"fc0880c2",
  1639 => x"fc0880ff",
  1640 => x"fffff806",
  1641 => x"555b7380",
  1642 => x"fffffff8",
  1643 => x"2e953880",
  1644 => x"c2fc08fe",
  1645 => x"0580ca88",
  1646 => x"082980ca",
  1647 => x"9c080557",
  1648 => x"b1c70480",
  1649 => x"547380c2",
  1650 => x"fc0c02b4",
  1651 => x"050d0402",
  1652 => x"f4050d74",
  1653 => x"70088105",
  1654 => x"710c7008",
  1655 => x"80ca8c08",
  1656 => x"06535371",
  1657 => x"8f388813",
  1658 => x"0851adfe",
  1659 => x"2d80c2fc",
  1660 => x"0888140c",
  1661 => x"810b80c2",
  1662 => x"fc0c028c",
  1663 => x"050d0402",
  1664 => x"f0050d75",
  1665 => x"881108fe",
  1666 => x"0580ca88",
  1667 => x"082980ca",
  1668 => x"9c081172",
  1669 => x"0880ca8c",
  1670 => x"08060579",
  1671 => x"55535454",
  1672 => x"a4ea2d02",
  1673 => x"90050d04",
  1674 => x"02f0050d",
  1675 => x"75881108",
  1676 => x"fe0580ca",
  1677 => x"88082980",
  1678 => x"ca9c0811",
  1679 => x"720880ca",
  1680 => x"8c080605",
  1681 => x"79555354",
  1682 => x"54a3a82d",
  1683 => x"0290050d",
  1684 => x"0402f405",
  1685 => x"0d747088",
  1686 => x"2a83fe80",
  1687 => x"06707298",
  1688 => x"2a077288",
  1689 => x"2b87fc80",
  1690 => x"80067398",
  1691 => x"2b81f00a",
  1692 => x"06717307",
  1693 => x"0780c2fc",
  1694 => x"0c565153",
  1695 => x"51028c05",
  1696 => x"0d0402f8",
  1697 => x"050d028e",
  1698 => x"0580f52d",
  1699 => x"74882b07",
  1700 => x"7083ffff",
  1701 => x"0680c2fc",
  1702 => x"0c510288",
  1703 => x"050d0402",
  1704 => x"f4050d74",
  1705 => x"76785354",
  1706 => x"52807125",
  1707 => x"97387270",
  1708 => x"81055480",
  1709 => x"f52d7270",
  1710 => x"81055481",
  1711 => x"b72dff11",
  1712 => x"5170eb38",
  1713 => x"807281b7",
  1714 => x"2d028c05",
  1715 => x"0d0402e8",
  1716 => x"050d7756",
  1717 => x"80705654",
  1718 => x"737624b6",
  1719 => x"3880ca94",
  1720 => x"08742eae",
  1721 => x"387351ae",
  1722 => x"f72d80c2",
  1723 => x"fc0880c2",
  1724 => x"fc080981",
  1725 => x"057080c2",
  1726 => x"fc08079f",
  1727 => x"2a770581",
  1728 => x"17575753",
  1729 => x"53747624",
  1730 => x"893880ca",
  1731 => x"94087426",
  1732 => x"d4387280",
  1733 => x"c2fc0c02",
  1734 => x"98050d04",
  1735 => x"02f0050d",
  1736 => x"80c2f808",
  1737 => x"1651b5ce",
  1738 => x"2d80c2fc",
  1739 => x"08802e9f",
  1740 => x"388b5380",
  1741 => x"c2fc0852",
  1742 => x"80c88451",
  1743 => x"b59f2d80",
  1744 => x"cac00854",
  1745 => x"73802e87",
  1746 => x"3880c884",
  1747 => x"51732d02",
  1748 => x"90050d04",
  1749 => x"02dc050d",
  1750 => x"80705a55",
  1751 => x"7480c2f8",
  1752 => x"0825b438",
  1753 => x"80ca9408",
  1754 => x"752eac38",
  1755 => x"7851aef7",
  1756 => x"2d80c2fc",
  1757 => x"08098105",
  1758 => x"7080c2fc",
  1759 => x"08079f2a",
  1760 => x"7605811b",
  1761 => x"5b565474",
  1762 => x"80c2f808",
  1763 => x"25893880",
  1764 => x"ca940879",
  1765 => x"26d63880",
  1766 => x"557880ca",
  1767 => x"94082781",
  1768 => x"db387851",
  1769 => x"aef72d80",
  1770 => x"c2fc0880",
  1771 => x"2e81ad38",
  1772 => x"80c2fc08",
  1773 => x"8b0580f5",
  1774 => x"2d70842a",
  1775 => x"70810677",
  1776 => x"1078842b",
  1777 => x"80c8840b",
  1778 => x"80f52d5c",
  1779 => x"5c535155",
  1780 => x"5673802e",
  1781 => x"80cb3874",
  1782 => x"16822bb9",
  1783 => x"a00b80c1",
  1784 => x"cc120c54",
  1785 => x"77753110",
  1786 => x"80cac411",
  1787 => x"55569074",
  1788 => x"70810556",
  1789 => x"81b72da0",
  1790 => x"7481b72d",
  1791 => x"7681ff06",
  1792 => x"81165854",
  1793 => x"73802e8a",
  1794 => x"389c5380",
  1795 => x"c88452b8",
  1796 => x"99048b53",
  1797 => x"80c2fc08",
  1798 => x"5280cac6",
  1799 => x"1651b8d4",
  1800 => x"04741682",
  1801 => x"2bb69c0b",
  1802 => x"80c1cc12",
  1803 => x"0c547681",
  1804 => x"ff068116",
  1805 => x"58547380",
  1806 => x"2e8a389c",
  1807 => x"5380c884",
  1808 => x"52b8cb04",
  1809 => x"8b5380c2",
  1810 => x"fc085277",
  1811 => x"75311080",
  1812 => x"cac40551",
  1813 => x"7655b59f",
  1814 => x"2db8f104",
  1815 => x"74902975",
  1816 => x"31701080",
  1817 => x"cac40551",
  1818 => x"5480c2fc",
  1819 => x"087481b7",
  1820 => x"2d811959",
  1821 => x"748b24a3",
  1822 => x"38b79904",
  1823 => x"74902975",
  1824 => x"31701080",
  1825 => x"cac4058c",
  1826 => x"77315751",
  1827 => x"54807481",
  1828 => x"b72d9e14",
  1829 => x"ff165654",
  1830 => x"74f33802",
  1831 => x"a4050d04",
  1832 => x"02fc050d",
  1833 => x"80c2f808",
  1834 => x"1351b5ce",
  1835 => x"2d80c2fc",
  1836 => x"08802e89",
  1837 => x"3880c2fc",
  1838 => x"0851a6cc",
  1839 => x"2d800b80",
  1840 => x"c2f80cb6",
  1841 => x"d42d92ad",
  1842 => x"2d028405",
  1843 => x"0d0402fc",
  1844 => x"050d7251",
  1845 => x"70fd2eb0",
  1846 => x"3870fd24",
  1847 => x"8a3870fc",
  1848 => x"2e80cc38",
  1849 => x"bab90470",
  1850 => x"fe2eb738",
  1851 => x"70ff2e09",
  1852 => x"810680c5",
  1853 => x"3880c2f8",
  1854 => x"08517080",
  1855 => x"2ebb38ff",
  1856 => x"1180c2f8",
  1857 => x"0cbab904",
  1858 => x"80c2f808",
  1859 => x"f0057080",
  1860 => x"c2f80c51",
  1861 => x"708025a1",
  1862 => x"38800b80",
  1863 => x"c2f80cba",
  1864 => x"b90480c2",
  1865 => x"f8088105",
  1866 => x"80c2f80c",
  1867 => x"bab90480",
  1868 => x"c2f80890",
  1869 => x"0580c2f8",
  1870 => x"0cb6d42d",
  1871 => x"92ad2d02",
  1872 => x"84050d04",
  1873 => x"02fc050d",
  1874 => x"800b80c2",
  1875 => x"f80cb6d4",
  1876 => x"2d91a92d",
  1877 => x"80c2fc08",
  1878 => x"80c2e80c",
  1879 => x"80c1c451",
  1880 => x"93d02d02",
  1881 => x"84050d04",
  1882 => x"7180cac0",
  1883 => x"0c040000",
  1884 => x"00ffffff",
  1885 => x"ff00ffff",
  1886 => x"ffff00ff",
  1887 => x"ffffff00",
  1888 => x"52657365",
  1889 => x"74204336",
  1890 => x"34000000",
  1891 => x"43363467",
  1892 => x"73206269",
  1893 => x"6f730000",
  1894 => x"41756469",
  1895 => x"6f206669",
  1896 => x"6c746572",
  1897 => x"00000000",
  1898 => x"4c6f6164",
  1899 => x"20443634",
  1900 => x"20646973",
  1901 => x"6b201000",
  1902 => x"44363420",
  1903 => x"72656164",
  1904 => x"206f6e6c",
  1905 => x"79000000",
  1906 => x"4c6f6164",
  1907 => x"20544150",
  1908 => x"20746170",
  1909 => x"65201000",
  1910 => x"45786974",
  1911 => x"00000000",
  1912 => x"48657820",
  1913 => x"64697370",
  1914 => x"2e207461",
  1915 => x"70652063",
  1916 => x"6f756e74",
  1917 => x"20757000",
  1918 => x"48657820",
  1919 => x"64697370",
  1920 => x"2e207461",
  1921 => x"70652063",
  1922 => x"6f756e74",
  1923 => x"20646f77",
  1924 => x"6e000000",
  1925 => x"48657820",
  1926 => x"64697370",
  1927 => x"2e206469",
  1928 => x"736b2074",
  1929 => x"7261636b",
  1930 => x"2d736563",
  1931 => x"746f7200",
  1932 => x"43494120",
  1933 => x"36323536",
  1934 => x"00000000",
  1935 => x"43494120",
  1936 => x"38353231",
  1937 => x"00000000",
  1938 => x"53494420",
  1939 => x"36353831",
  1940 => x"204d6f6e",
  1941 => x"6f000000",
  1942 => x"53494420",
  1943 => x"36353831",
  1944 => x"20537465",
  1945 => x"72656f00",
  1946 => x"53494420",
  1947 => x"38353830",
  1948 => x"204d6f6e",
  1949 => x"6f000000",
  1950 => x"53494420",
  1951 => x"38353830",
  1952 => x"20537465",
  1953 => x"72656f00",
  1954 => x"53494420",
  1955 => x"50736575",
  1956 => x"646f2053",
  1957 => x"74657265",
  1958 => x"6f000000",
  1959 => x"524f4d20",
  1960 => x"6c6f6164",
  1961 => x"696e6720",
  1962 => x"6661696c",
  1963 => x"65640000",
  1964 => x"4f4b0000",
  1965 => x"496e6974",
  1966 => x"69616c69",
  1967 => x"7a696e67",
  1968 => x"20534420",
  1969 => x"63617264",
  1970 => x"0a000000",
  1971 => x"16200000",
  1972 => x"14200000",
  1973 => x"15200000",
  1974 => x"53442069",
  1975 => x"6e69742e",
  1976 => x"2e2e0a00",
  1977 => x"53442063",
  1978 => x"61726420",
  1979 => x"72657365",
  1980 => x"74206661",
  1981 => x"696c6564",
  1982 => x"210a0000",
  1983 => x"53444843",
  1984 => x"20657272",
  1985 => x"6f72210a",
  1986 => x"00000000",
  1987 => x"57726974",
  1988 => x"65206661",
  1989 => x"696c6564",
  1990 => x"0a000000",
  1991 => x"52656164",
  1992 => x"20666169",
  1993 => x"6c65640a",
  1994 => x"00000000",
  1995 => x"43617264",
  1996 => x"20696e69",
  1997 => x"74206661",
  1998 => x"696c6564",
  1999 => x"0a000000",
  2000 => x"46415431",
  2001 => x"36202020",
  2002 => x"00000000",
  2003 => x"46415433",
  2004 => x"32202020",
  2005 => x"00000000",
  2006 => x"4e6f2070",
  2007 => x"61727469",
  2008 => x"74696f6e",
  2009 => x"20736967",
  2010 => x"0a000000",
  2011 => x"42616420",
  2012 => x"70617274",
  2013 => x"0a000000",
  2014 => x"4261636b",
  2015 => x"00000000",
  2016 => x"00000002",
  2017 => x"ffffffff",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000002",
  2025 => x"00001d80",
  2026 => x"00000304",
  2027 => x"00000001",
  2028 => x"00001d8c",
  2029 => x"00000000",
  2030 => x"00000003",
  2031 => x"00002038",
  2032 => x"00000005",
  2033 => x"00000001",
  2034 => x"00001d98",
  2035 => x"00000001",
  2036 => x"00000003",
  2037 => x"00002030",
  2038 => x"00000002",
  2039 => x"00000002",
  2040 => x"00001da8",
  2041 => x"0000031b",
  2042 => x"00000001",
  2043 => x"00001db8",
  2044 => x"00000002",
  2045 => x"00000002",
  2046 => x"00001dc8",
  2047 => x"0000032e",
  2048 => x"00000003",
  2049 => x"00002024",
  2050 => x"00000003",
  2051 => x"00000002",
  2052 => x"00001dd8",
  2053 => x"000008c6",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00001de0",
  2058 => x"00001df8",
  2059 => x"00001e14",
  2060 => x"00001e30",
  2061 => x"00001e3c",
  2062 => x"00001e48",
  2063 => x"00001e58",
  2064 => x"00001e68",
  2065 => x"00001e78",
  2066 => x"00001e88",
  2067 => x"00000004",
  2068 => x"00001e9c",
  2069 => x"0000204c",
  2070 => x"00000004",
  2071 => x"00001eb0",
  2072 => x"00001fa0",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000002",
  2098 => x"00002544",
  2099 => x"00001b1c",
  2100 => x"00000002",
  2101 => x"00002562",
  2102 => x"00001b1c",
  2103 => x"00000002",
  2104 => x"00002580",
  2105 => x"00001b1c",
  2106 => x"00000002",
  2107 => x"0000259e",
  2108 => x"00001b1c",
  2109 => x"00000002",
  2110 => x"000025bc",
  2111 => x"00001b1c",
  2112 => x"00000002",
  2113 => x"000025da",
  2114 => x"00001b1c",
  2115 => x"00000002",
  2116 => x"000025f8",
  2117 => x"00001b1c",
  2118 => x"00000002",
  2119 => x"00002616",
  2120 => x"00001b1c",
  2121 => x"00000002",
  2122 => x"00002634",
  2123 => x"00001b1c",
  2124 => x"00000002",
  2125 => x"00002652",
  2126 => x"00001b1c",
  2127 => x"00000002",
  2128 => x"00002670",
  2129 => x"00001b1c",
  2130 => x"00000002",
  2131 => x"0000268e",
  2132 => x"00001b1c",
  2133 => x"00000002",
  2134 => x"000026ac",
  2135 => x"00001b1c",
  2136 => x"00000004",
  2137 => x"00001f78",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00001cce",
  2142 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

